
`include "../Design/wrt_controller.v"
`include "../Design/rd_controller.v"
module design_top #(parameter N=32)(
     
     input m_axi_lite_aclk,                 //IP to master
     input m_axi_lite_aresetn,              //active low reset IP to master

     //READ OPERATION WITHOUT ERROR
 
//---------------------------------IP to Master -------------------------------------------------
//
//
     input IP2Bus_MstRd_Req,                 //read request from IP to Master
     input [N-1:0]IP2Bus_Mst_rAddr,           //address for both read and write IP to master
     
     input [N-1:0]IP2Bus_Mst_wrAddr,           //address for both read and write IP to master
                    //   For Write operations   //
     
     input [N-1:0]IP2Bus_MstWr_d,
     input IP2Bus_MstWr_Req,
     input [(N/8)-1:0]IP2Bus_Mst_BE,

//----------------------------------------------------------------------------------------------
//
//
//---------------------------------Master to Slave --------------------------------------------- 

     output [N-1:0]m_axi_lite_araddr,        //address--> ouput from master to slave
     output m_axi_lite_arvalid,              //valid signal generate by master to slave
     output m_axi_lite_rready,               // ready signal generated by master to slave for reading data from slave

                    //   For Write operations   //

     output [N-1:0]m_axi_lite_awaddr,
     output [2:0]m_axi_lite_awprot,
     output m_axi_lite_awvalid,
     output [N-1:0]m_axi_lite_wdata,
     output [(N/8)-1:0]m_axi_lite_wstrb,
     output m_axi_lite_wvalid,
     output m_axi_lite_bready,
//----------------------------------------------------------------------------------------------
//
//
//--------------------------------- Slave to Master --------------------------------------------- 
     
     input m_axi_lite_arready,               //ip==> Ready signal generated from slave to master
     input [N-1:0]m_axi_lite_rdata,          //ip==> data generated from particular address from slave to master
     input m_axi_lite_rvalid,                // valid signal from slave to master for transferring data 
    // utput i
     input [1:0]m_axi_lite_resp,             //from slave to master to known that was operation OK or not

                    //   For Write operations   //


     input m_axi_lite_awready,
     input m_axi_lite_wready,
     input [1:0]m_axi_lite_bresp,
     input m_axi_lite_bvalid,

//----------------------------------------------------------------------------------------------
//
//
//--------------------------------- Master to IP --------------------------------------------- 

     output [N-1:0]Bus2IP_MstRd_d,      //output from master to IP containing Data
     output Bus2IP_Mst_wrCmdAck,        //acknowledge signal from master to IP after succesfully reading address
     output Bus2IP_Mst_wrCmplt,         //From Master to IP , When data is fetched
     
     output Bus2IP_Mst_rCmdAck,         //acknowledge signal from master to IP after succesfully reading address
     output Bus2IP_Mst_rCmplt,        //From Master to IP , When data is fetched

     output Bus2IP_Mst_Src_Rdy_n,    //Active low,generated from master to IP,indicating data asserted on bus is valid
     output BUS2IP_Mstwr_Dst_Rdy_n,  //Active low,generated from master to IP,indicating data asserted on bus is valid
     output md_error,                 //Active high master detected error output discrete. 
     output BUS2IP_Mst_rError,

     output BUS2IP_Mst_wrError);
//----------------------------------------------------------------------------------------------
  assign md_error = md_error_r | md_error_w;
rd_controller rdc(


///--------------------------------- Master to IP --------------------------------------------- 

     Bus2IP_MstRd_d,           //output from master to IP containing Data
     Bus2IP_Mst_rCmdAck,               //acknowledge signal from master to IP after succesfully reading address
     Bus2IP_Mst_rCmplt,                //From Master to IP , When data is fetched

     Bus2IP_Mst_Src_Rdy_n,            //Active low , generated from master to IP,indicating data asserted on bus is valid
     md_error_r,                        //Active high master detected error output discrete. 
     BUS2IP_Mst_rError,
//----------------------------------------------------------------------------------------------
//
//
//---------------------------------Master to Slave --------------------------------------------- 
 
     m_axi_lite_araddr,        //address--> ouput from master to slave
     m_axi_lite_arvalid,              //valid signal generate by master to slave
     m_axi_lite_rready,               // ready signal generated by master to slave for reading data from slave

//----------------------------------------------------------------------------------------------
//
//
//---------------------------------IP to Master -------------------------------------------------

     m_axi_lite_aclk,                  //IP to master
     m_axi_lite_aresetn,               //active low reset IP to master
     
     IP2Bus_MstRd_Req,                 //read request from IP to Master
     IP2Bus_Mst_rAddr,           //address for both read and write IP to master
     
//----------------------------------------------------------------------------------------------
//
//
//--------------------------------- Slave to Master --------------------------------------------- 
     
     m_axi_lite_arready,               //ip==> Ready signal generated from slave to master
     m_axi_lite_rdata,          //ip==> data generated from particular address from slave to master
     m_axi_lite_rvalid,                // valid signal from slave to master for transferring data 
     m_axi_lite_resp             //from slave to master to known that was operation OK or not

//----------------------------------------------------------------------------------------------
//
);


wrt_controller wrc(
                        

//MAster to Slave
     m_axi_lite_awaddr, //address--> ouput from master to slave
     m_axi_lite_awvalid, //valid signal generate by master to slave
     m_axi_lite_wdata, //data --> master to slave--through IP
     m_axi_lite_wvalid, // valid signal generated by master to slave for writing data from slave
     m_axi_lite_wstrb, //strobe from master to slave --> through IP
     m_axi_lite_bready, //ready signal from master to slave -- for getting response signal


// Master to IP

     Bus2IP_Mst_wrCmdAck, //acknowledge signal from master to IP after succesfully reading address
     Bus2IP_Mst_wrCmplt, //From Master to IP , When data is fetched
     Bus2IP_Mst_dst_Rdy_n, //Active low , generated from master to IP,indicating data asserted on bus is valid
     md_error_w, //Active high master detected error output discrete 
     BUS2IP_Mst_wrError, 


     m_axi_lite_aclk, //IP to master
     m_axi_lite_aresetn, //active low reset IP to master
 
//IP to Master
     IP2Bus_MstWr_Req, //write request from IP to Master
     IP2Bus_Mst_wrAddr, //address for both read and write IP to master
     IP2Bus_MstWr_d, //write data from ip to bus
     IP2Bus_Mst_BE, // strobe signal from ip to bus

//Slave to Master
     m_axi_lite_awready, //ip==> Ready signal generated to get data from  master
     m_axi_lite_wready, //ip==> ready signal generated to get data from master
     m_axi_lite_bvalid, // valid response signal from slave to master for transferring response signal to master 
     m_axi_lite_bresp   //from slave to master to known that was operation OK or not
     );






endmodule
