  module rd_controller #(parameter N=32)(

///--------------------------------- Master to IP --------------------------------------------- 
     output reg [N-1:0]Bus2IP_MstRd_d,           //output from master to IP containing Data
     output reg Bus2IP_Mst_CmdAck,               //acknowledge signal from master to IP after succesfully reading address
     output reg Bus2IP_Mst_Cmplt,                //From Master to IP , When data is fetched
     output reg Bus2IP_Mst_Src_Rdy_n,            //Active low , generated from master to IP,indicating data asserted on bus is valid
     output reg md_error,                        //Active high master detected error output discrete. 
     output reg BUS2IP_Mst_Error,
//----------------------------------------------------------------------------------------------
//
//
//---------------------------------Master to Slave --------------------------------------------- 

     output reg [N-1:0]m_axi_lite_araddr,        //address--> ouput from master to slave
     output reg m_axi_lite_arvalid,              //valid signal generate by master to slave
     output reg m_axi_lite_rready,               // ready signal generated by master to slave for reading data from slave

//----------------------------------------------------------------------------------------------
//
//
//---------------------------------IP to Master -------------------------------------------------

     input m_axi_lite_aclk,                  //IP to master
     input m_axi_lite_aresetn,               //active low reset IP to master
     input IP2Bus_MstRd_Req,                 //read request from IP to Master
     input [N-1:0]IP2Bus_Mst_Addr,           //address for both read and write IP to master
     
//----------------------------------------------------------------------------------------------
//
//
//--------------------------------- Slave to Master --------------------------------------------- 
     
     input m_axi_lite_arready,               //ip==> Ready signal generated from slave to master
     input [N-1:0]m_axi_lite_rdata,          //ip==> data generated from particular address from slave to master
     input m_axi_lite_rvalid,                // valid signal from slave to master for transferring data 
     input [1:0]m_axi_lite_resp             //from slave to master to known that was operation OK or not

//----------------------------------------------------------------------------------------------
//
);

     reg [1:0] next_state,present_state;  //  State variables that required for moore state machine
     parameter s0 = 2'b00;
     parameter s1 = 2'b01;
     parameter s2 = 2'b10;
     parameter s3 = 2'b11;

     always @(posedge m_axi_lite_aclk, negedge m_axi_lite_aresetn) begin
          if (!m_axi_lite_aresetn)
            next_state=s0;
          else 
            present_state=next_state;

          case (present_state) 
               s0:  begin
                    //$display("I'm in state 0");
                    if (IP2Bus_MstRd_Req)
                         next_state=s1;
                    else if(m_axi_lite_aresetn)
                         next_state=s0;
               end

               s1:  begin
                    //$display("I'm in state 1");
                    if (m_axi_lite_arready)  begin
                         m_axi_lite_araddr = IP2Bus_Mst_Addr;
                         next_state = s2;
                    end
               end

               s2:  begin
                    //$display("I'm in state 2");
                    if (m_axi_lite_rvalid)   begin
                         next_state = s3;
                    end
               end

               s3:  begin
                    //$display("I'm in state 3");
                    next_state = s0;
               end                            
          endcase
     end


     always @(present_state) begin
          case(present_state)   
               s0:  begin                 
                    Bus2IP_MstRd_d <= 0;           //output from master to IP containing Data
                    Bus2IP_Mst_CmdAck<=0;               //acknowledge signal from master to IP after succesfully reading address
                    Bus2IP_Mst_Cmplt<=0;                //From Master to IP , When data is fetched

                    Bus2IP_Mst_Src_Rdy_n<=1;            //Active low , generated from master to IP,indicating data asserted on bus is valid
                    md_error<=0;                        //Active high master detected error output discrete. 

                    //m_axi_lite_araddr <= 0;        //address--> ouput from master to slave
                    m_axi_lite_arvalid <= 0;              //valid signal generate by master to slave
                    m_axi_lite_rready <= 0;               // ready signal generated by master to slave for reading data from slave
               end

               s1:  begin
                    m_axi_lite_rready<=1;
                    m_axi_lite_arvalid<=1;
               end

               s2:  begin
                    m_axi_lite_arvalid<=0;
                    Bus2IP_Mst_CmdAck<=1;
                    @(posedge m_axi_lite_aclk) ;
                    Bus2IP_Mst_CmdAck<= 0;
               end

               s3:  begin
                    Bus2IP_Mst_CmdAck<=0;
                    if (m_axi_lite_resp>0) begin
                         md_error<=1;
                         BUS2IP_Mst_Error<=1;
                    end
                    Bus2IP_Mst_Cmplt<=1;
                    Bus2IP_MstRd_d <=  m_axi_lite_rdata;
                    Bus2IP_Mst_Src_Rdy_n <= 0;

               end
          endcase  
     end          
     endmodule
